
`timescale 1ns / 1ps
module Sine_LUT ( step, val );
	input [9:0] step;
	output reg [9:0] val;
	always @ (step) begin
		case (step)
			10'd0: val <= 10'd1023;
			10'd1: val <= 10'd1029;
			10'd2: val <= 10'd1036;
			10'd3: val <= 10'd1042;
			10'd4: val <= 10'd1048;
			10'd5: val <= 10'd1054;
			10'd6: val <= 10'd1061;
			10'd7: val <= 10'd1067;
			10'd8: val <= 10'd1073;
			10'd9: val <= 10'd1079;
			10'd10: val <= 10'd1086;
			10'd11: val <= 10'd1092;
			10'd12: val <= 10'd1098;
			10'd13: val <= 10'd1105;
			10'd14: val <= 10'd1111;
			10'd15: val <= 10'd1117;
			10'd16: val <= 10'd1123;
			10'd17: val <= 10'd1130;
			10'd18: val <= 10'd1136;
			10'd19: val <= 10'd1142;
			10'd20: val <= 10'd1148;
			10'd21: val <= 10'd1154;
			10'd22: val <= 10'd1161;
			10'd23: val <= 10'd1167;
			10'd24: val <= 10'd1173;
			10'd25: val <= 10'd1179;
			10'd26: val <= 10'd1186;
			10'd27: val <= 10'd1192;
			10'd28: val <= 10'd1198;
			10'd29: val <= 10'd1204;
			10'd30: val <= 10'd1210;
			10'd31: val <= 10'd1216;
			10'd32: val <= 10'd1223;
			10'd33: val <= 10'd1229;
			10'd34: val <= 10'd1235;
			10'd35: val <= 10'd1241;
			10'd36: val <= 10'd1247;
			10'd37: val <= 10'd1253;
			10'd38: val <= 10'd1259;
			10'd39: val <= 10'd1265;
			10'd40: val <= 10'd1272;
			10'd41: val <= 10'd1278;
			10'd42: val <= 10'd1284;
			10'd43: val <= 10'd1290;
			10'd44: val <= 10'd1296;
			10'd45: val <= 10'd1302;
			10'd46: val <= 10'd1308;
			10'd47: val <= 10'd1314;
			10'd48: val <= 10'd1320;
			10'd49: val <= 10'd1326;
			10'd50: val <= 10'd1332;
			10'd51: val <= 10'd1338;
			10'd52: val <= 10'd1344;
			10'd53: val <= 10'd1350;
			10'd54: val <= 10'd1356;
			10'd55: val <= 10'd1362;
			10'd56: val <= 10'd1368;
			10'd57: val <= 10'd1374;
			10'd58: val <= 10'd1379;
			10'd59: val <= 10'd1385;
			10'd60: val <= 10'd1391;
			10'd61: val <= 10'd1397;
			10'd62: val <= 10'd1403;
			10'd63: val <= 10'd1409;
			10'd64: val <= 10'd1414;
			10'd65: val <= 10'd1420;
			10'd66: val <= 10'd1426;
			10'd67: val <= 10'd1432;
			10'd68: val <= 10'd1438;
			10'd69: val <= 10'd1443;
			10'd70: val <= 10'd1449;
			10'd71: val <= 10'd1455;
			10'd72: val <= 10'd1460;
			10'd73: val <= 10'd1466;
			10'd74: val <= 10'd1472;
			10'd75: val <= 10'd1477;
			10'd76: val <= 10'd1483;
			10'd77: val <= 10'd1489;
			10'd78: val <= 10'd1494;
			10'd79: val <= 10'd1500;
			10'd80: val <= 10'd1505;
			10'd81: val <= 10'd1511;
			10'd82: val <= 10'd1516;
			10'd83: val <= 10'd1522;
			10'd84: val <= 10'd1527;
			10'd85: val <= 10'd1533;
			10'd86: val <= 10'd1538;
			10'd87: val <= 10'd1544;
			10'd88: val <= 10'd1549;
			10'd89: val <= 10'd1554;
			10'd90: val <= 10'd1560;
			10'd91: val <= 10'd1565;
			10'd92: val <= 10'd1570;
			10'd93: val <= 10'd1576;
			10'd94: val <= 10'd1581;
			10'd95: val <= 10'd1586;
			10'd96: val <= 10'd1591;
			10'd97: val <= 10'd1597;
			10'd98: val <= 10'd1602;
			10'd99: val <= 10'd1607;
			10'd100: val <= 10'd1612;
			10'd101: val <= 10'd1617;
			10'd102: val <= 10'd1622;
			10'd103: val <= 10'd1627;
			10'd104: val <= 10'd1632;
			10'd105: val <= 10'd1637;
			10'd106: val <= 10'd1642;
			10'd107: val <= 10'd1647;
			10'd108: val <= 10'd1652;
			10'd109: val <= 10'd1657;
			10'd110: val <= 10'd1662;
			10'd111: val <= 10'd1667;
			10'd112: val <= 10'd1672;
			10'd113: val <= 10'd1677;
			10'd114: val <= 10'd1682;
			10'd115: val <= 10'd1686;
			10'd116: val <= 10'd1691;
			10'd117: val <= 10'd1696;
			10'd118: val <= 10'd1701;
			10'd119: val <= 10'd1705;
			10'd120: val <= 10'd1710;
			10'd121: val <= 10'd1715;
			10'd122: val <= 10'd1719;
			10'd123: val <= 10'd1724;
			10'd124: val <= 10'd1728;
			10'd125: val <= 10'd1733;
			10'd126: val <= 10'd1737;
			10'd127: val <= 10'd1742;
			10'd128: val <= 10'd1746;
			10'd129: val <= 10'd1751;
			10'd130: val <= 10'd1755;
			10'd131: val <= 10'd1760;
			10'd132: val <= 10'd1764;
			10'd133: val <= 10'd1768;
			10'd134: val <= 10'd1773;
			10'd135: val <= 10'd1777;
			10'd136: val <= 10'd1781;
			10'd137: val <= 10'd1785;
			10'd138: val <= 10'd1789;
			10'd139: val <= 10'd1794;
			10'd140: val <= 10'd1798;
			10'd141: val <= 10'd1802;
			10'd142: val <= 10'd1806;
			10'd143: val <= 10'd1810;
			10'd144: val <= 10'd1814;
			10'd145: val <= 10'd1818;
			10'd146: val <= 10'd1822;
			10'd147: val <= 10'd1826;
			10'd148: val <= 10'd1829;
			10'd149: val <= 10'd1833;
			10'd150: val <= 10'd1837;
			10'd151: val <= 10'd1841;
			10'd152: val <= 10'd1845;
			10'd153: val <= 10'd1848;
			10'd154: val <= 10'd1852;
			10'd155: val <= 10'd1856;
			10'd156: val <= 10'd1859;
			10'd157: val <= 10'd1863;
			10'd158: val <= 10'd1867;
			10'd159: val <= 10'd1870;
			10'd160: val <= 10'd1874;
			10'd161: val <= 10'd1877;
			10'd162: val <= 10'd1881;
			10'd163: val <= 10'd1884;
			10'd164: val <= 10'd1887;
			10'd165: val <= 10'd1891;
			10'd166: val <= 10'd1894;
			10'd167: val <= 10'd1897;
			10'd168: val <= 10'd1900;
			10'd169: val <= 10'd1904;
			10'd170: val <= 10'd1907;
			10'd171: val <= 10'd1910;
			10'd172: val <= 10'd1913;
			10'd173: val <= 10'd1916;
			10'd174: val <= 10'd1919;
			10'd175: val <= 10'd1922;
			10'd176: val <= 10'd1925;
			10'd177: val <= 10'd1928;
			10'd178: val <= 10'd1931;
			10'd179: val <= 10'd1934;
			10'd180: val <= 10'd1937;
			10'd181: val <= 10'd1940;
			10'd182: val <= 10'd1942;
			10'd183: val <= 10'd1945;
			10'd184: val <= 10'd1948;
			10'd185: val <= 10'd1950;
			10'd186: val <= 10'd1953;
			10'd187: val <= 10'd1956;
			10'd188: val <= 10'd1958;
			10'd189: val <= 10'd1961;
			10'd190: val <= 10'd1963;
			10'd191: val <= 10'd1966;
			10'd192: val <= 10'd1968;
			10'd193: val <= 10'd1971;
			10'd194: val <= 10'd1973;
			10'd195: val <= 10'd1975;
			10'd196: val <= 10'd1977;
			10'd197: val <= 10'd1980;
			10'd198: val <= 10'd1982;
			10'd199: val <= 10'd1984;
			10'd200: val <= 10'd1986;
			10'd201: val <= 10'd1988;
			10'd202: val <= 10'd1990;
			10'd203: val <= 10'd1992;
			10'd204: val <= 10'd1994;
			10'd205: val <= 10'd1996;
			10'd206: val <= 10'd1998;
			10'd207: val <= 10'd2000;
			10'd208: val <= 10'd2002;
			10'd209: val <= 10'd2004;
			10'd210: val <= 10'd2006;
			10'd211: val <= 10'd2007;
			10'd212: val <= 10'd2009;
			10'd213: val <= 10'd2011;
			10'd214: val <= 10'd2012;
			10'd215: val <= 10'd2014;
			10'd216: val <= 10'd2015;
			10'd217: val <= 10'd2017;
			10'd218: val <= 10'd2018;
			10'd219: val <= 10'd2020;
			10'd220: val <= 10'd2021;
			10'd221: val <= 10'd2022;
			10'd222: val <= 10'd2024;
			10'd223: val <= 10'd2025;
			10'd224: val <= 10'd2026;
			10'd225: val <= 10'd2028;
			10'd226: val <= 10'd2029;
			10'd227: val <= 10'd2030;
			10'd228: val <= 10'd2031;
			10'd229: val <= 10'd2032;
			10'd230: val <= 10'd2033;
			10'd231: val <= 10'd2034;
			10'd232: val <= 10'd2035;
			10'd233: val <= 10'd2036;
			10'd234: val <= 10'd2037;
			10'd235: val <= 10'd2038;
			10'd236: val <= 10'd2038;
			10'd237: val <= 10'd2039;
			10'd238: val <= 10'd2040;
			10'd239: val <= 10'd2040;
			10'd240: val <= 10'd2041;
			10'd241: val <= 10'd2042;
			10'd242: val <= 10'd2042;
			10'd243: val <= 10'd2043;
			10'd244: val <= 10'd2043;
			10'd245: val <= 10'd2044;
			10'd246: val <= 10'd2044;
			10'd247: val <= 10'd2044;
			10'd248: val <= 10'd2045;
			10'd249: val <= 10'd2045;
			10'd250: val <= 10'd2045;
			10'd251: val <= 10'd2046;
			10'd252: val <= 10'd2046;
			10'd253: val <= 10'd2046;
			10'd254: val <= 10'd2046;
			10'd255: val <= 10'd2046;
			10'd256: val <= 10'd2046;
			10'd257: val <= 10'd2046;
			10'd258: val <= 10'd2046;
			10'd259: val <= 10'd2046;
			10'd260: val <= 10'd2046;
			10'd261: val <= 10'd2046;
			10'd262: val <= 10'd2045;
			10'd263: val <= 10'd2045;
			10'd264: val <= 10'd2045;
			10'd265: val <= 10'd2044;
			10'd266: val <= 10'd2044;
			10'd267: val <= 10'd2044;
			10'd268: val <= 10'd2043;
			10'd269: val <= 10'd2043;
			10'd270: val <= 10'd2042;
			10'd271: val <= 10'd2042;
			10'd272: val <= 10'd2041;
			10'd273: val <= 10'd2040;
			10'd274: val <= 10'd2040;
			10'd275: val <= 10'd2039;
			10'd276: val <= 10'd2038;
			10'd277: val <= 10'd2038;
			10'd278: val <= 10'd2037;
			10'd279: val <= 10'd2036;
			10'd280: val <= 10'd2035;
			10'd281: val <= 10'd2034;
			10'd282: val <= 10'd2033;
			10'd283: val <= 10'd2032;
			10'd284: val <= 10'd2031;
			10'd285: val <= 10'd2030;
			10'd286: val <= 10'd2029;
			10'd287: val <= 10'd2028;
			10'd288: val <= 10'd2026;
			10'd289: val <= 10'd2025;
			10'd290: val <= 10'd2024;
			10'd291: val <= 10'd2022;
			10'd292: val <= 10'd2021;
			10'd293: val <= 10'd2020;
			10'd294: val <= 10'd2018;
			10'd295: val <= 10'd2017;
			10'd296: val <= 10'd2015;
			10'd297: val <= 10'd2014;
			10'd298: val <= 10'd2012;
			10'd299: val <= 10'd2011;
			10'd300: val <= 10'd2009;
			10'd301: val <= 10'd2007;
			10'd302: val <= 10'd2006;
			10'd303: val <= 10'd2004;
			10'd304: val <= 10'd2002;
			10'd305: val <= 10'd2000;
			10'd306: val <= 10'd1998;
			10'd307: val <= 10'd1996;
			10'd308: val <= 10'd1994;
			10'd309: val <= 10'd1992;
			10'd310: val <= 10'd1990;
			10'd311: val <= 10'd1988;
			10'd312: val <= 10'd1986;
			10'd313: val <= 10'd1984;
			10'd314: val <= 10'd1982;
			10'd315: val <= 10'd1980;
			10'd316: val <= 10'd1977;
			10'd317: val <= 10'd1975;
			10'd318: val <= 10'd1973;
			10'd319: val <= 10'd1971;
			10'd320: val <= 10'd1968;
			10'd321: val <= 10'd1966;
			10'd322: val <= 10'd1963;
			10'd323: val <= 10'd1961;
			10'd324: val <= 10'd1958;
			10'd325: val <= 10'd1956;
			10'd326: val <= 10'd1953;
			10'd327: val <= 10'd1950;
			10'd328: val <= 10'd1948;
			10'd329: val <= 10'd1945;
			10'd330: val <= 10'd1942;
			10'd331: val <= 10'd1940;
			10'd332: val <= 10'd1937;
			10'd333: val <= 10'd1934;
			10'd334: val <= 10'd1931;
			10'd335: val <= 10'd1928;
			10'd336: val <= 10'd1925;
			10'd337: val <= 10'd1922;
			10'd338: val <= 10'd1919;
			10'd339: val <= 10'd1916;
			10'd340: val <= 10'd1913;
			10'd341: val <= 10'd1910;
			10'd342: val <= 10'd1907;
			10'd343: val <= 10'd1904;
			10'd344: val <= 10'd1900;
			10'd345: val <= 10'd1897;
			10'd346: val <= 10'd1894;
			10'd347: val <= 10'd1891;
			10'd348: val <= 10'd1887;
			10'd349: val <= 10'd1884;
			10'd350: val <= 10'd1881;
			10'd351: val <= 10'd1877;
			10'd352: val <= 10'd1874;
			10'd353: val <= 10'd1870;
			10'd354: val <= 10'd1867;
			10'd355: val <= 10'd1863;
			10'd356: val <= 10'd1859;
			10'd357: val <= 10'd1856;
			10'd358: val <= 10'd1852;
			10'd359: val <= 10'd1848;
			10'd360: val <= 10'd1845;
			10'd361: val <= 10'd1841;
			10'd362: val <= 10'd1837;
			10'd363: val <= 10'd1833;
			10'd364: val <= 10'd1829;
			10'd365: val <= 10'd1826;
			10'd366: val <= 10'd1822;
			10'd367: val <= 10'd1818;
			10'd368: val <= 10'd1814;
			10'd369: val <= 10'd1810;
			10'd370: val <= 10'd1806;
			10'd371: val <= 10'd1802;
			10'd372: val <= 10'd1798;
			10'd373: val <= 10'd1794;
			10'd374: val <= 10'd1789;
			10'd375: val <= 10'd1785;
			10'd376: val <= 10'd1781;
			10'd377: val <= 10'd1777;
			10'd378: val <= 10'd1773;
			10'd379: val <= 10'd1768;
			10'd380: val <= 10'd1764;
			10'd381: val <= 10'd1760;
			10'd382: val <= 10'd1755;
			10'd383: val <= 10'd1751;
			10'd384: val <= 10'd1746;
			10'd385: val <= 10'd1742;
			10'd386: val <= 10'd1737;
			10'd387: val <= 10'd1733;
			10'd388: val <= 10'd1728;
			10'd389: val <= 10'd1724;
			10'd390: val <= 10'd1719;
			10'd391: val <= 10'd1715;
			10'd392: val <= 10'd1710;
			10'd393: val <= 10'd1705;
			10'd394: val <= 10'd1701;
			10'd395: val <= 10'd1696;
			10'd396: val <= 10'd1691;
			10'd397: val <= 10'd1686;
			10'd398: val <= 10'd1682;
			10'd399: val <= 10'd1677;
			10'd400: val <= 10'd1672;
			10'd401: val <= 10'd1667;
			10'd402: val <= 10'd1662;
			10'd403: val <= 10'd1657;
			10'd404: val <= 10'd1652;
			10'd405: val <= 10'd1647;
			10'd406: val <= 10'd1642;
			10'd407: val <= 10'd1637;
			10'd408: val <= 10'd1632;
			10'd409: val <= 10'd1627;
			10'd410: val <= 10'd1622;
			10'd411: val <= 10'd1617;
			10'd412: val <= 10'd1612;
			10'd413: val <= 10'd1607;
			10'd414: val <= 10'd1602;
			10'd415: val <= 10'd1597;
			10'd416: val <= 10'd1591;
			10'd417: val <= 10'd1586;
			10'd418: val <= 10'd1581;
			10'd419: val <= 10'd1576;
			10'd420: val <= 10'd1570;
			10'd421: val <= 10'd1565;
			10'd422: val <= 10'd1560;
			10'd423: val <= 10'd1554;
			10'd424: val <= 10'd1549;
			10'd425: val <= 10'd1544;
			10'd426: val <= 10'd1538;
			10'd427: val <= 10'd1533;
			10'd428: val <= 10'd1527;
			10'd429: val <= 10'd1522;
			10'd430: val <= 10'd1516;
			10'd431: val <= 10'd1511;
			10'd432: val <= 10'd1505;
			10'd433: val <= 10'd1500;
			10'd434: val <= 10'd1494;
			10'd435: val <= 10'd1489;
			10'd436: val <= 10'd1483;
			10'd437: val <= 10'd1477;
			10'd438: val <= 10'd1472;
			10'd439: val <= 10'd1466;
			10'd440: val <= 10'd1460;
			10'd441: val <= 10'd1455;
			10'd442: val <= 10'd1449;
			10'd443: val <= 10'd1443;
			10'd444: val <= 10'd1438;
			10'd445: val <= 10'd1432;
			10'd446: val <= 10'd1426;
			10'd447: val <= 10'd1420;
			10'd448: val <= 10'd1414;
			10'd449: val <= 10'd1409;
			10'd450: val <= 10'd1403;
			10'd451: val <= 10'd1397;
			10'd452: val <= 10'd1391;
			10'd453: val <= 10'd1385;
			10'd454: val <= 10'd1379;
			10'd455: val <= 10'd1374;
			10'd456: val <= 10'd1368;
			10'd457: val <= 10'd1362;
			10'd458: val <= 10'd1356;
			10'd459: val <= 10'd1350;
			10'd460: val <= 10'd1344;
			10'd461: val <= 10'd1338;
			10'd462: val <= 10'd1332;
			10'd463: val <= 10'd1326;
			10'd464: val <= 10'd1320;
			10'd465: val <= 10'd1314;
			10'd466: val <= 10'd1308;
			10'd467: val <= 10'd1302;
			10'd468: val <= 10'd1296;
			10'd469: val <= 10'd1290;
			10'd470: val <= 10'd1284;
			10'd471: val <= 10'd1278;
			10'd472: val <= 10'd1272;
			10'd473: val <= 10'd1265;
			10'd474: val <= 10'd1259;
			10'd475: val <= 10'd1253;
			10'd476: val <= 10'd1247;
			10'd477: val <= 10'd1241;
			10'd478: val <= 10'd1235;
			10'd479: val <= 10'd1229;
			10'd480: val <= 10'd1223;
			10'd481: val <= 10'd1216;
			10'd482: val <= 10'd1210;
			10'd483: val <= 10'd1204;
			10'd484: val <= 10'd1198;
			10'd485: val <= 10'd1192;
			10'd486: val <= 10'd1186;
			10'd487: val <= 10'd1179;
			10'd488: val <= 10'd1173;
			10'd489: val <= 10'd1167;
			10'd490: val <= 10'd1161;
			10'd491: val <= 10'd1154;
			10'd492: val <= 10'd1148;
			10'd493: val <= 10'd1142;
			10'd494: val <= 10'd1136;
			10'd495: val <= 10'd1130;
			10'd496: val <= 10'd1123;
			10'd497: val <= 10'd1117;
			10'd498: val <= 10'd1111;
			10'd499: val <= 10'd1105;
			10'd500: val <= 10'd1098;
			10'd501: val <= 10'd1092;
			10'd502: val <= 10'd1086;
			10'd503: val <= 10'd1079;
			10'd504: val <= 10'd1073;
			10'd505: val <= 10'd1067;
			10'd506: val <= 10'd1061;
			10'd507: val <= 10'd1054;
			10'd508: val <= 10'd1048;
			10'd509: val <= 10'd1042;
			10'd510: val <= 10'd1036;
			10'd511: val <= 10'd1029;
			10'd512: val <= 10'd1023;
			10'd513: val <= 10'd1017;
			10'd514: val <= 10'd1010;
			10'd515: val <= 10'd1004;
			10'd516: val <= 10'd998;
			10'd517: val <= 10'd992;
			10'd518: val <= 10'd985;
			10'd519: val <= 10'd979;
			10'd520: val <= 10'd973;
			10'd521: val <= 10'd967;
			10'd522: val <= 10'd960;
			10'd523: val <= 10'd954;
			10'd524: val <= 10'd948;
			10'd525: val <= 10'd941;
			10'd526: val <= 10'd935;
			10'd527: val <= 10'd929;
			10'd528: val <= 10'd923;
			10'd529: val <= 10'd916;
			10'd530: val <= 10'd910;
			10'd531: val <= 10'd904;
			10'd532: val <= 10'd898;
			10'd533: val <= 10'd892;
			10'd534: val <= 10'd885;
			10'd535: val <= 10'd879;
			10'd536: val <= 10'd873;
			10'd537: val <= 10'd867;
			10'd538: val <= 10'd860;
			10'd539: val <= 10'd854;
			10'd540: val <= 10'd848;
			10'd541: val <= 10'd842;
			10'd542: val <= 10'd836;
			10'd543: val <= 10'd830;
			10'd544: val <= 10'd823;
			10'd545: val <= 10'd817;
			10'd546: val <= 10'd811;
			10'd547: val <= 10'd805;
			10'd548: val <= 10'd799;
			10'd549: val <= 10'd793;
			10'd550: val <= 10'd787;
			10'd551: val <= 10'd781;
			10'd552: val <= 10'd774;
			10'd553: val <= 10'd768;
			10'd554: val <= 10'd762;
			10'd555: val <= 10'd756;
			10'd556: val <= 10'd750;
			10'd557: val <= 10'd744;
			10'd558: val <= 10'd738;
			10'd559: val <= 10'd732;
			10'd560: val <= 10'd726;
			10'd561: val <= 10'd720;
			10'd562: val <= 10'd714;
			10'd563: val <= 10'd708;
			10'd564: val <= 10'd702;
			10'd565: val <= 10'd696;
			10'd566: val <= 10'd690;
			10'd567: val <= 10'd684;
			10'd568: val <= 10'd678;
			10'd569: val <= 10'd672;
			10'd570: val <= 10'd667;
			10'd571: val <= 10'd661;
			10'd572: val <= 10'd655;
			10'd573: val <= 10'd649;
			10'd574: val <= 10'd643;
			10'd575: val <= 10'd637;
			10'd576: val <= 10'd632;
			10'd577: val <= 10'd626;
			10'd578: val <= 10'd620;
			10'd579: val <= 10'd614;
			10'd580: val <= 10'd608;
			10'd581: val <= 10'd603;
			10'd582: val <= 10'd597;
			10'd583: val <= 10'd591;
			10'd584: val <= 10'd586;
			10'd585: val <= 10'd580;
			10'd586: val <= 10'd574;
			10'd587: val <= 10'd569;
			10'd588: val <= 10'd563;
			10'd589: val <= 10'd557;
			10'd590: val <= 10'd552;
			10'd591: val <= 10'd546;
			10'd592: val <= 10'd541;
			10'd593: val <= 10'd535;
			10'd594: val <= 10'd530;
			10'd595: val <= 10'd524;
			10'd596: val <= 10'd519;
			10'd597: val <= 10'd513;
			10'd598: val <= 10'd508;
			10'd599: val <= 10'd502;
			10'd600: val <= 10'd497;
			10'd601: val <= 10'd492;
			10'd602: val <= 10'd486;
			10'd603: val <= 10'd481;
			10'd604: val <= 10'd476;
			10'd605: val <= 10'd470;
			10'd606: val <= 10'd465;
			10'd607: val <= 10'd460;
			10'd608: val <= 10'd455;
			10'd609: val <= 10'd449;
			10'd610: val <= 10'd444;
			10'd611: val <= 10'd439;
			10'd612: val <= 10'd434;
			10'd613: val <= 10'd429;
			10'd614: val <= 10'd424;
			10'd615: val <= 10'd419;
			10'd616: val <= 10'd414;
			10'd617: val <= 10'd409;
			10'd618: val <= 10'd404;
			10'd619: val <= 10'd399;
			10'd620: val <= 10'd394;
			10'd621: val <= 10'd389;
			10'd622: val <= 10'd384;
			10'd623: val <= 10'd379;
			10'd624: val <= 10'd374;
			10'd625: val <= 10'd369;
			10'd626: val <= 10'd364;
			10'd627: val <= 10'd360;
			10'd628: val <= 10'd355;
			10'd629: val <= 10'd350;
			10'd630: val <= 10'd345;
			10'd631: val <= 10'd341;
			10'd632: val <= 10'd336;
			10'd633: val <= 10'd331;
			10'd634: val <= 10'd327;
			10'd635: val <= 10'd322;
			10'd636: val <= 10'd318;
			10'd637: val <= 10'd313;
			10'd638: val <= 10'd309;
			10'd639: val <= 10'd304;
			10'd640: val <= 10'd300;
			10'd641: val <= 10'd295;
			10'd642: val <= 10'd291;
			10'd643: val <= 10'd286;
			10'd644: val <= 10'd282;
			10'd645: val <= 10'd278;
			10'd646: val <= 10'd273;
			10'd647: val <= 10'd269;
			10'd648: val <= 10'd265;
			10'd649: val <= 10'd261;
			10'd650: val <= 10'd257;
			10'd651: val <= 10'd252;
			10'd652: val <= 10'd248;
			10'd653: val <= 10'd244;
			10'd654: val <= 10'd240;
			10'd655: val <= 10'd236;
			10'd656: val <= 10'd232;
			10'd657: val <= 10'd228;
			10'd658: val <= 10'd224;
			10'd659: val <= 10'd220;
			10'd660: val <= 10'd217;
			10'd661: val <= 10'd213;
			10'd662: val <= 10'd209;
			10'd663: val <= 10'd205;
			10'd664: val <= 10'd201;
			10'd665: val <= 10'd198;
			10'd666: val <= 10'd194;
			10'd667: val <= 10'd190;
			10'd668: val <= 10'd187;
			10'd669: val <= 10'd183;
			10'd670: val <= 10'd179;
			10'd671: val <= 10'd176;
			10'd672: val <= 10'd172;
			10'd673: val <= 10'd169;
			10'd674: val <= 10'd165;
			10'd675: val <= 10'd162;
			10'd676: val <= 10'd159;
			10'd677: val <= 10'd155;
			10'd678: val <= 10'd152;
			10'd679: val <= 10'd149;
			10'd680: val <= 10'd146;
			10'd681: val <= 10'd142;
			10'd682: val <= 10'd139;
			10'd683: val <= 10'd136;
			10'd684: val <= 10'd133;
			10'd685: val <= 10'd130;
			10'd686: val <= 10'd127;
			10'd687: val <= 10'd124;
			10'd688: val <= 10'd121;
			10'd689: val <= 10'd118;
			10'd690: val <= 10'd115;
			10'd691: val <= 10'd112;
			10'd692: val <= 10'd109;
			10'd693: val <= 10'd106;
			10'd694: val <= 10'd104;
			10'd695: val <= 10'd101;
			10'd696: val <= 10'd98;
			10'd697: val <= 10'd96;
			10'd698: val <= 10'd93;
			10'd699: val <= 10'd90;
			10'd700: val <= 10'd88;
			10'd701: val <= 10'd85;
			10'd702: val <= 10'd83;
			10'd703: val <= 10'd80;
			10'd704: val <= 10'd78;
			10'd705: val <= 10'd75;
			10'd706: val <= 10'd73;
			10'd707: val <= 10'd71;
			10'd708: val <= 10'd69;
			10'd709: val <= 10'd66;
			10'd710: val <= 10'd64;
			10'd711: val <= 10'd62;
			10'd712: val <= 10'd60;
			10'd713: val <= 10'd58;
			10'd714: val <= 10'd56;
			10'd715: val <= 10'd54;
			10'd716: val <= 10'd52;
			10'd717: val <= 10'd50;
			10'd718: val <= 10'd48;
			10'd719: val <= 10'd46;
			10'd720: val <= 10'd44;
			10'd721: val <= 10'd42;
			10'd722: val <= 10'd40;
			10'd723: val <= 10'd39;
			10'd724: val <= 10'd37;
			10'd725: val <= 10'd35;
			10'd726: val <= 10'd34;
			10'd727: val <= 10'd32;
			10'd728: val <= 10'd31;
			10'd729: val <= 10'd29;
			10'd730: val <= 10'd28;
			10'd731: val <= 10'd26;
			10'd732: val <= 10'd25;
			10'd733: val <= 10'd24;
			10'd734: val <= 10'd22;
			10'd735: val <= 10'd21;
			10'd736: val <= 10'd20;
			10'd737: val <= 10'd18;
			10'd738: val <= 10'd17;
			10'd739: val <= 10'd16;
			10'd740: val <= 10'd15;
			10'd741: val <= 10'd14;
			10'd742: val <= 10'd13;
			10'd743: val <= 10'd12;
			10'd744: val <= 10'd11;
			10'd745: val <= 10'd10;
			10'd746: val <= 10'd9;
			10'd747: val <= 10'd8;
			10'd748: val <= 10'd8;
			10'd749: val <= 10'd7;
			10'd750: val <= 10'd6;
			10'd751: val <= 10'd6;
			10'd752: val <= 10'd5;
			10'd753: val <= 10'd4;
			10'd754: val <= 10'd4;
			10'd755: val <= 10'd3;
			10'd756: val <= 10'd3;
			10'd757: val <= 10'd2;
			10'd758: val <= 10'd2;
			10'd759: val <= 10'd2;
			10'd760: val <= 10'd1;
			10'd761: val <= 10'd1;
			10'd762: val <= 10'd1;
			10'd763: val <= 10'd0;
			10'd764: val <= 10'd0;
			10'd765: val <= 10'd0;
			10'd766: val <= 10'd0;
			10'd767: val <= 10'd0;
			10'd768: val <= 10'd0;
			10'd769: val <= 10'd0;
			10'd770: val <= 10'd0;
			10'd771: val <= 10'd0;
			10'd772: val <= 10'd0;
			10'd773: val <= 10'd0;
			10'd774: val <= 10'd1;
			10'd775: val <= 10'd1;
			10'd776: val <= 10'd1;
			10'd777: val <= 10'd2;
			10'd778: val <= 10'd2;
			10'd779: val <= 10'd2;
			10'd780: val <= 10'd3;
			10'd781: val <= 10'd3;
			10'd782: val <= 10'd4;
			10'd783: val <= 10'd4;
			10'd784: val <= 10'd5;
			10'd785: val <= 10'd6;
			10'd786: val <= 10'd6;
			10'd787: val <= 10'd7;
			10'd788: val <= 10'd8;
			10'd789: val <= 10'd8;
			10'd790: val <= 10'd9;
			10'd791: val <= 10'd10;
			10'd792: val <= 10'd11;
			10'd793: val <= 10'd12;
			10'd794: val <= 10'd13;
			10'd795: val <= 10'd14;
			10'd796: val <= 10'd15;
			10'd797: val <= 10'd16;
			10'd798: val <= 10'd17;
			10'd799: val <= 10'd18;
			10'd800: val <= 10'd20;
			10'd801: val <= 10'd21;
			10'd802: val <= 10'd22;
			10'd803: val <= 10'd24;
			10'd804: val <= 10'd25;
			10'd805: val <= 10'd26;
			10'd806: val <= 10'd28;
			10'd807: val <= 10'd29;
			10'd808: val <= 10'd31;
			10'd809: val <= 10'd32;
			10'd810: val <= 10'd34;
			10'd811: val <= 10'd35;
			10'd812: val <= 10'd37;
			10'd813: val <= 10'd39;
			10'd814: val <= 10'd40;
			10'd815: val <= 10'd42;
			10'd816: val <= 10'd44;
			10'd817: val <= 10'd46;
			10'd818: val <= 10'd48;
			10'd819: val <= 10'd50;
			10'd820: val <= 10'd52;
			10'd821: val <= 10'd54;
			10'd822: val <= 10'd56;
			10'd823: val <= 10'd58;
			10'd824: val <= 10'd60;
			10'd825: val <= 10'd62;
			10'd826: val <= 10'd64;
			10'd827: val <= 10'd66;
			10'd828: val <= 10'd69;
			10'd829: val <= 10'd71;
			10'd830: val <= 10'd73;
			10'd831: val <= 10'd75;
			10'd832: val <= 10'd78;
			10'd833: val <= 10'd80;
			10'd834: val <= 10'd83;
			10'd835: val <= 10'd85;
			10'd836: val <= 10'd88;
			10'd837: val <= 10'd90;
			10'd838: val <= 10'd93;
			10'd839: val <= 10'd96;
			10'd840: val <= 10'd98;
			10'd841: val <= 10'd101;
			10'd842: val <= 10'd104;
			10'd843: val <= 10'd106;
			10'd844: val <= 10'd109;
			10'd845: val <= 10'd112;
			10'd846: val <= 10'd115;
			10'd847: val <= 10'd118;
			10'd848: val <= 10'd121;
			10'd849: val <= 10'd124;
			10'd850: val <= 10'd127;
			10'd851: val <= 10'd130;
			10'd852: val <= 10'd133;
			10'd853: val <= 10'd136;
			10'd854: val <= 10'd139;
			10'd855: val <= 10'd142;
			10'd856: val <= 10'd146;
			10'd857: val <= 10'd149;
			10'd858: val <= 10'd152;
			10'd859: val <= 10'd155;
			10'd860: val <= 10'd159;
			10'd861: val <= 10'd162;
			10'd862: val <= 10'd165;
			10'd863: val <= 10'd169;
			10'd864: val <= 10'd172;
			10'd865: val <= 10'd176;
			10'd866: val <= 10'd179;
			10'd867: val <= 10'd183;
			10'd868: val <= 10'd187;
			10'd869: val <= 10'd190;
			10'd870: val <= 10'd194;
			10'd871: val <= 10'd198;
			10'd872: val <= 10'd201;
			10'd873: val <= 10'd205;
			10'd874: val <= 10'd209;
			10'd875: val <= 10'd213;
			10'd876: val <= 10'd217;
			10'd877: val <= 10'd220;
			10'd878: val <= 10'd224;
			10'd879: val <= 10'd228;
			10'd880: val <= 10'd232;
			10'd881: val <= 10'd236;
			10'd882: val <= 10'd240;
			10'd883: val <= 10'd244;
			10'd884: val <= 10'd248;
			10'd885: val <= 10'd252;
			10'd886: val <= 10'd257;
			10'd887: val <= 10'd261;
			10'd888: val <= 10'd265;
			10'd889: val <= 10'd269;
			10'd890: val <= 10'd273;
			10'd891: val <= 10'd278;
			10'd892: val <= 10'd282;
			10'd893: val <= 10'd286;
			10'd894: val <= 10'd291;
			10'd895: val <= 10'd295;
			10'd896: val <= 10'd300;
			10'd897: val <= 10'd304;
			10'd898: val <= 10'd309;
			10'd899: val <= 10'd313;
			10'd900: val <= 10'd318;
			10'd901: val <= 10'd322;
			10'd902: val <= 10'd327;
			10'd903: val <= 10'd331;
			10'd904: val <= 10'd336;
			10'd905: val <= 10'd341;
			10'd906: val <= 10'd345;
			10'd907: val <= 10'd350;
			10'd908: val <= 10'd355;
			10'd909: val <= 10'd360;
			10'd910: val <= 10'd364;
			10'd911: val <= 10'd369;
			10'd912: val <= 10'd374;
			10'd913: val <= 10'd379;
			10'd914: val <= 10'd384;
			10'd915: val <= 10'd389;
			10'd916: val <= 10'd394;
			10'd917: val <= 10'd399;
			10'd918: val <= 10'd404;
			10'd919: val <= 10'd409;
			10'd920: val <= 10'd414;
			10'd921: val <= 10'd419;
			10'd922: val <= 10'd424;
			10'd923: val <= 10'd429;
			10'd924: val <= 10'd434;
			10'd925: val <= 10'd439;
			10'd926: val <= 10'd444;
			10'd927: val <= 10'd449;
			10'd928: val <= 10'd455;
			10'd929: val <= 10'd460;
			10'd930: val <= 10'd465;
			10'd931: val <= 10'd470;
			10'd932: val <= 10'd476;
			10'd933: val <= 10'd481;
			10'd934: val <= 10'd486;
			10'd935: val <= 10'd492;
			10'd936: val <= 10'd497;
			10'd937: val <= 10'd502;
			10'd938: val <= 10'd508;
			10'd939: val <= 10'd513;
			10'd940: val <= 10'd519;
			10'd941: val <= 10'd524;
			10'd942: val <= 10'd530;
			10'd943: val <= 10'd535;
			10'd944: val <= 10'd541;
			10'd945: val <= 10'd546;
			10'd946: val <= 10'd552;
			10'd947: val <= 10'd557;
			10'd948: val <= 10'd563;
			10'd949: val <= 10'd569;
			10'd950: val <= 10'd574;
			10'd951: val <= 10'd580;
			10'd952: val <= 10'd586;
			10'd953: val <= 10'd591;
			10'd954: val <= 10'd597;
			10'd955: val <= 10'd603;
			10'd956: val <= 10'd608;
			10'd957: val <= 10'd614;
			10'd958: val <= 10'd620;
			10'd959: val <= 10'd626;
			10'd960: val <= 10'd632;
			10'd961: val <= 10'd637;
			10'd962: val <= 10'd643;
			10'd963: val <= 10'd649;
			10'd964: val <= 10'd655;
			10'd965: val <= 10'd661;
			10'd966: val <= 10'd667;
			10'd967: val <= 10'd672;
			10'd968: val <= 10'd678;
			10'd969: val <= 10'd684;
			10'd970: val <= 10'd690;
			10'd971: val <= 10'd696;
			10'd972: val <= 10'd702;
			10'd973: val <= 10'd708;
			10'd974: val <= 10'd714;
			10'd975: val <= 10'd720;
			10'd976: val <= 10'd726;
			10'd977: val <= 10'd732;
			10'd978: val <= 10'd738;
			10'd979: val <= 10'd744;
			10'd980: val <= 10'd750;
			10'd981: val <= 10'd756;
			10'd982: val <= 10'd762;
			10'd983: val <= 10'd768;
			10'd984: val <= 10'd774;
			10'd985: val <= 10'd781;
			10'd986: val <= 10'd787;
			10'd987: val <= 10'd793;
			10'd988: val <= 10'd799;
			10'd989: val <= 10'd805;
			10'd990: val <= 10'd811;
			10'd991: val <= 10'd817;
			10'd992: val <= 10'd823;
			10'd993: val <= 10'd830;
			10'd994: val <= 10'd836;
			10'd995: val <= 10'd842;
			10'd996: val <= 10'd848;
			10'd997: val <= 10'd854;
			10'd998: val <= 10'd860;
			10'd999: val <= 10'd867;
			10'd1000: val <= 10'd873;
			10'd1001: val <= 10'd879;
			10'd1002: val <= 10'd885;
			10'd1003: val <= 10'd892;
			10'd1004: val <= 10'd898;
			10'd1005: val <= 10'd904;
			10'd1006: val <= 10'd910;
			10'd1007: val <= 10'd916;
			10'd1008: val <= 10'd923;
			10'd1009: val <= 10'd929;
			10'd1010: val <= 10'd935;
			10'd1011: val <= 10'd941;
			10'd1012: val <= 10'd948;
			10'd1013: val <= 10'd954;
			10'd1014: val <= 10'd960;
			10'd1015: val <= 10'd967;
			10'd1016: val <= 10'd973;
			10'd1017: val <= 10'd979;
			10'd1018: val <= 10'd985;
			10'd1019: val <= 10'd992;
			10'd1020: val <= 10'd998;
			10'd1021: val <= 10'd1004;
			10'd1022: val <= 10'd1010;
			10'd1023: val <= 10'd1017;
		endcase
	end
endmodule

module Sine_LUT_TEST ( );
	reg [10:0] step;
	wire [10:0] val;
	Sine_LUT UUT (step, val);
	initial begin
		$dumpvars;
		step <= 0;
		#100
		repeat (9) begin
			#10 step <= step + 1;
		end
	end
endmodule